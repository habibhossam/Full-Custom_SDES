* SPICE NETLIST
***************************************

.SUBCKT GND
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT VDD
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT Inverter_1 Vdd Gnd Out In
** N=4 EP=4 IP=3 FDC=2
M0 Out In Gnd Gnd NMOS25 L=2.5e-07 W=7.5e-07 AD=4.875e-13 AS=4.875e-13 PD=2.8e-06 PS=2.8e-06 $X=205 $Y=-1630 $D=1
M1 Out In Vdd Vdd PMOS25 L=2.5e-07 W=1.5e-06 AD=9.75e-13 AS=9.75e-13 PD=4.3e-06 PS=4.3e-06 $X=205 $Y=855 $D=2
.ENDS
***************************************
.SUBCKT pmos25x_Auto_6_1
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B S D G
.ENDS
***************************************
.SUBCKT nmos25x_Auto_5_1
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: S D B G
.ENDS
***************************************
.SUBCKT XOR Vdd Out Gnd A B
** N=11 EP=5 IP=44 FDC=12
M0 6 10 Out Gnd NMOS25 L=2.5e-07 W=1.5e-06 AD=5.625e-13 AS=9.75e-13 PD=2.25e-06 PS=4.3e-06 $X=7105 $Y=-775 $D=1
M1 Gnd 11 6 Gnd NMOS25 L=2.5e-07 W=1.5e-06 AD=5.625e-13 AS=5.625e-13 PD=2.25e-06 PS=2.25e-06 $X=8105 $Y=-775 $D=1
M2 7 B Gnd Gnd NMOS25 L=2.5e-07 W=1.5e-06 AD=5.625e-13 AS=5.625e-13 PD=2.25e-06 PS=2.25e-06 $X=9105 $Y=-775 $D=1
M3 Out A 7 Gnd NMOS25 L=2.5e-07 W=1.5e-06 AD=9.75e-13 AS=5.625e-13 PD=4.3e-06 PS=2.25e-06 $X=10105 $Y=-775 $D=1
M4 8 A Vdd Vdd PMOS25 L=2.5e-07 W=3e-06 AD=1.125e-12 AS=1.95e-12 PD=3.75e-06 PS=7.3e-06 $X=7105 $Y=10320 $D=2
M5 Out 11 8 Vdd PMOS25 L=2.5e-07 W=3e-06 AD=1.125e-12 AS=1.125e-12 PD=3.75e-06 PS=3.75e-06 $X=8105 $Y=10320 $D=2
M6 9 B Out Vdd PMOS25 L=2.5e-07 W=3e-06 AD=1.125e-12 AS=1.125e-12 PD=3.75e-06 PS=3.75e-06 $X=9105 $Y=10320 $D=2
M7 Vdd 10 9 Vdd PMOS25 L=2.5e-07 W=3e-06 AD=1.95e-12 AS=1.125e-12 PD=7.3e-06 PS=3.75e-06 $X=10105 $Y=10320 $D=2
X8 Vdd Gnd 11 B Inverter_1 $T=905 2320 0 0 $X=-2085 $Y=-995
X9 Vdd Gnd 10 A Inverter_1 $T=905 11435 0 0 $X=-2085 $Y=8120
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6 7 8
*.CALIBRE ICV_CELL 9
** N=8 EP=8 IP=10 FDC=24
X0 3 4 1 7 2 XOR $T=0 0 0 0 $X=-5000 $Y=-4855
X1 3 6 1 8 5 XOR $T=0 21280 0 0 $X=-5000 $Y=16425
.ENDS
***************************************
.SUBCKT pmos25x_Auto_7_1 B S D G
** N=5 EP=4 IP=0 FDC=1
M0 D G S B PMOS25 L=2.5e-07 W=1.5e-06 AD=5.625e-13 AS=9.75e-13 PD=2.25e-06 PS=4.3e-06 $X=0 $Y=0 $D=2
.ENDS
***************************************
.SUBCKT nand_2 Vdd Gnd Out A B
** N=6 EP=5 IP=21 FDC=4
M0 6 A Gnd Gnd NMOS25 L=2.5e-07 W=1.5e-06 AD=5.625e-13 AS=9.75e-13 PD=2.25e-06 PS=4.3e-06 $X=705 $Y=-1355 $D=1
M1 Out B 6 Gnd NMOS25 L=2.5e-07 W=1.5e-06 AD=9.75e-13 AS=5.625e-13 PD=4.3e-06 PS=2.25e-06 $X=1705 $Y=-1355 $D=1
X6 Vdd Vdd Out A pmos25x_Auto_7_1 $T=705 2630 0 0 $X=-695 $Y=1880
X7 Vdd Vdd Out B pmos25x_Auto_7_1 $T=1955 2630 1 180 $X=305 $Y=1880
.ENDS
***************************************
.SUBCKT pmos25x_Auto_8_1
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: B S D G
.ENDS
***************************************
.SUBCKT nmos25x_Auto_9_1 S D B G
** N=4 EP=4 IP=0 FDC=1
M0 D G S B NMOS25 L=2.5e-07 W=7.5e-07 AD=2.8125e-13 AS=4.875e-13 PD=1.5e-06 PS=2.8e-06 $X=0 $Y=0 $D=1
.ENDS
***************************************
.SUBCKT nor_2 Vdd Out Gnd A B
** N=6 EP=5 IP=18 FDC=4
M0 6 A Vdd Vdd PMOS25 L=2.5e-07 W=1.5e-06 AD=5.625e-13 AS=9.75e-13 PD=2.25e-06 PS=4.3e-06 $X=4505 $Y=3955 $D=2
M1 Out B 6 Vdd PMOS25 L=2.5e-07 W=1.5e-06 AD=9.75e-13 AS=5.625e-13 PD=4.3e-06 PS=2.25e-06 $X=5505 $Y=3955 $D=2
X4 Gnd Out Gnd A nmos25x_Auto_9_1 $T=4505 820 0 0 $X=3605 $Y=-480
X5 Gnd Out Gnd B nmos25x_Auto_9_1 $T=5755 820 1 180 $X=4605 $Y=-480
.ENDS
***************************************
.SUBCKT AND_2 Gnd A B Vdd Y
** N=6 EP=5 IP=9 FDC=6
X0 Vdd Gnd Y 6 Inverter_1 $T=8800 3840 0 0 $X=5810 $Y=525
X1 Vdd Gnd 6 A B nand_2 $T=0 2295 0 0 $X=-1475 $Y=-1745
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7
*.CALIBRE ICV_CELL 9
** N=7 EP=7 IP=10 FDC=12
X0 1 3 4 2 5 AND_2 $T=0 0 0 0 $X=-1475 $Y=-1745
X1 1 5 6 2 7 AND_2 $T=13370 0 0 0 $X=11895 $Y=-1745
.ENDS
***************************************
.SUBCKT S1 Gnd Vdd I3 I0 I2 I1 S11 S10
** N=35 EP=8 IP=114 FDC=134
X0 Vdd Gnd 9 I3 Inverter_1 $T=21045 2945 0 0 $X=18055 $Y=-370
X1 Vdd Gnd 10 I3 Inverter_1 $T=21045 136020 1 0 $X=18055 $Y=131530
X2 Vdd Gnd 11 I0 Inverter_1 $T=26595 2945 0 0 $X=23605 $Y=-370
X3 Vdd Gnd 12 I0 Inverter_1 $T=26595 136020 1 0 $X=23605 $Y=131530
X4 Vdd Gnd 13 I2 Inverter_1 $T=32150 2945 0 0 $X=29160 $Y=-370
X5 Vdd Gnd 14 I1 Inverter_1 $T=32150 136020 1 0 $X=29160 $Y=131530
X6 Vdd Gnd 15 I1 Inverter_1 $T=37680 2945 0 0 $X=34690 $Y=-370
X7 Vdd Gnd S11 30 33 nand_2 $T=73635 86330 1 0 $X=72160 $Y=79015
X8 Vdd Gnd S10 34 35 nand_2 $T=79470 51740 0 0 $X=77995 $Y=47700
X9 Vdd 30 Gnd 25 29 nor_2 $T=62790 87565 1 0 $X=65895 $Y=80310
X10 Vdd 33 Gnd 24 28 nor_2 $T=62790 111320 1 0 $X=65895 $Y=104065
X11 Vdd 35 Gnd 26 31 nor_2 $T=68625 26750 0 0 $X=71730 $Y=26270
X12 Vdd 34 Gnd 27 32 nor_2 $T=68625 50505 0 0 $X=71730 $Y=50025
X13 Gnd Vdd I1 10 16 12 25 ICV_2 $T=38590 88250 1 0 $X=37115 $Y=78640
X14 Gnd Vdd I0 10 17 I2 29 ICV_2 $T=38590 100105 1 0 $X=37115 $Y=90495
X15 Gnd Vdd I0 I3 18 I1 24 ICV_2 $T=38590 111960 1 0 $X=37115 $Y=102350
X16 Gnd Vdd 14 I3 19 12 28 ICV_2 $T=38590 123815 1 0 $X=37115 $Y=114205
X17 Gnd Vdd 15 I3 20 13 31 ICV_2 $T=44455 14250 0 0 $X=42980 $Y=12505
X18 Gnd Vdd I0 I2 21 I1 26 ICV_2 $T=44455 26105 0 0 $X=42980 $Y=24360
X19 Gnd Vdd I0 13 22 15 32 ICV_2 $T=44455 37960 0 0 $X=42980 $Y=36215
X20 Gnd Vdd I2 9 23 11 27 ICV_2 $T=44455 49815 0 0 $X=42980 $Y=48070
.ENDS
***************************************
.SUBCKT ICV_3 1 2 3 4 5 6 7 8 9 10 11
*.CALIBRE ICV_CELL 9
** N=11 EP=11 IP=14 FDC=24
X0 1 2 3 4 5 6 7 ICV_2 $T=0 0 0 0 $X=-1475 $Y=-1745
X1 1 2 3 8 9 10 11 ICV_2 $T=0 11855 0 0 $X=-1475 $Y=10110
.ENDS
***************************************
.SUBCKT S00 Gnd Vdd A B C D S0_0
** N=25 EP=7 IP=69 FDC=86
X0 Vdd Gnd 8 A Inverter_1 $T=6555 -9080 0 0 $X=3565 $Y=-12395
X1 Vdd Gnd 9 B Inverter_1 $T=12105 -9080 0 0 $X=9115 $Y=-12395
X2 Vdd Gnd 10 C Inverter_1 $T=17660 -9080 0 0 $X=14670 $Y=-12395
X3 Vdd Gnd 11 D Inverter_1 $T=23190 -9080 0 0 $X=20200 $Y=-12395
X4 Vdd Gnd 22 21 Inverter_1 $T=72330 27130 0 0 $X=69340 $Y=23815
X5 Vdd Gnd S0_0 23 24 nand_2 $T=74445 49505 0 0 $X=72970 $Y=45465
X6 Vdd 21 Gnd 17 19 nor_2 $T=58480 24365 0 0 $X=61585 $Y=23885
X7 Vdd 23 Gnd 18 20 nor_2 $T=59915 48095 0 0 $X=63020 $Y=47615
X8 Vdd 24 Gnd 22 25 nor_2 $T=76150 24330 0 0 $X=79255 $Y=23850
X9 Gnd Vdd A B 16 11 18 ICV_2 $T=32950 47420 0 0 $X=31475 $Y=45675
X10 Gnd Vdd 8 9 12 C 25 B 13 10 19 ICV_3 $T=32950 0 0 0 $X=31475 $Y=-1745
X11 Gnd Vdd A 9 14 D 17 C 15 D 20 ICV_3 $T=32950 23710 0 0 $X=31475 $Y=21965
.ENDS
***************************************
.SUBCKT ICV_4 1 2 3 4 5
*.CALIBRE ICV_CELL 9
** N=5 EP=5 IP=8 FDC=4
X0 2 1 3 5 Inverter_1 $T=0 0 0 0 $X=-2990 $Y=-3315
X1 2 1 4 3 Inverter_1 $T=5155 0 0 0 $X=2165 $Y=-3315
.ENDS
***************************************
.SUBCKT FK Gnd k7 k6 k5 k4 I7 I6 I5 I4 I3 I2 I1 I0 k0 k1 k2 Vdd O3 O2 O1
+ O0 k3 23 24 O4 O5 O6 O7
** N=54 EP=28 IP=146 FDC=436
X0 Vdd Gnd 41 40 Inverter_1 $T=23578 157710 0 0 $X=20588 $Y=154395
X1 Vdd Gnd 42 37 Inverter_1 $T=29128 157710 0 0 $X=26138 $Y=154395
X2 Vdd Gnd 43 39 Inverter_1 $T=34683 157710 0 0 $X=31693 $Y=154395
X3 Vdd Gnd 44 38 Inverter_1 $T=40213 157710 0 0 $X=37223 $Y=154395
X4 Vdd O5 Gnd I5 24 XOR $T=106835 156910 0 0 $X=101835 $Y=152055
X5 Vdd O4 Gnd I4 54 XOR $T=106855 178190 0 0 $X=101855 $Y=173335
X6 Gnd I0 Vdd 40 I3 39 k7 k6 ICV_1 $T=-3750 71790 0 0 $X=-8750 $Y=66935
X7 Gnd I2 Vdd 38 I1 37 k5 k4 ICV_1 $T=-3750 114350 0 0 $X=-8750 $Y=109495
X8 Gnd I2 Vdd 36 I1 35 k3 k2 ICV_1 $T=-3750 156910 0 0 $X=-8750 $Y=152055
X9 Gnd I0 Vdd 34 I3 33 k1 k0 ICV_1 $T=-3750 199470 0 0 $X=-8750 $Y=194615
X10 Gnd 53 Vdd O7 23 O6 I7 I6 ICV_1 $T=106835 114350 0 0 $X=101835 $Y=109495
X11 Vdd Gnd 53 51 52 nand_2 $T=85958 210735 0 0 $X=84483 $Y=206695
X12 Vdd 52 Gnd 47 50 nor_2 $T=71513 185215 0 0 $X=74618 $Y=184735
X13 Vdd 51 Gnd 48 49 nor_2 $T=71513 208985 0 0 $X=74618 $Y=208505
X14 Gnd 44 39 Vdd 50 AND_2 $T=48863 172815 0 0 $X=47388 $Y=171070
X15 Gnd 40 42 Vdd 45 AND_2 $T=48863 184670 0 0 $X=47388 $Y=182925
X16 Gnd 41 44 Vdd 49 AND_2 $T=48863 196525 0 0 $X=47388 $Y=194780
X17 Gnd 40 37 Vdd 46 AND_2 $T=48863 208380 0 0 $X=47388 $Y=206635
X18 Gnd 45 39 Vdd 47 AND_2 $T=62233 184670 0 0 $X=60758 $Y=182925
X19 Gnd 46 43 Vdd 48 AND_2 $T=62233 208380 0 0 $X=60758 $Y=206635
X20 Gnd Vdd 36 33 35 34 23 24 S1 $T=6415 11080 0 0 $X=24470 $Y=10710
X21 Gnd Vdd 40 37 39 38 54 S00 $T=17023 280510 1 0 $X=20528 $Y=220595
X22 Gnd Vdd 29 O1 I1 ICV_4 $T=-18830 187890 0 0 $X=-21820 $Y=184575
X23 Gnd Vdd 30 O0 I0 ICV_4 $T=-18830 206405 0 0 $X=-21820 $Y=203090
X24 Gnd Vdd 31 O2 I2 ICV_4 $T=-18815 163880 0 0 $X=-21805 $Y=160565
X25 Gnd Vdd 32 O3 I3 ICV_4 $T=-18815 232515 0 0 $X=-21805 $Y=229200
.ENDS
***************************************
.SUBCKT SDES Gnd K1 K3 K6 K2 K7 K0 K4 K9 I6 I7 I0 I4 I2 I5 I3 I1 Vdd K5 K8
+ O7 O5 O2 O6 O1 O4 O0 O3
** N=40 EP=28 IP=56 FDC=872
X0 Gnd K9 K3 K1 K6 I6 I2 I5 I7 I4 I0 I3 I1 K4 K0 K7 Vdd 28 27 26
+ 25 K2 19 20 21 22 23 24
+ FK $T=-13843 27130 0 0 $X=-57295 $Y=31820
X1 Gnd K2 K7 K4 K5 28 27 26 25 24 23 22 21 K9 K1 K8 Vdd O4 O0 O3
+ O1 K0 31 32 O7 O5 O2 O6
+ FK $T=189540 27130 0 0 $X=146088 $Y=31820
.ENDS
***************************************
